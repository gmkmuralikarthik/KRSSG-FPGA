// Verilog test fixture created from schematic /home/ise/ism_projects/xi share/KRSSG FPGA CODES/cordic_test/test.sch - Sat Feb 29 04:25:32 2020

`timescale 1ns / 1ps

module test_test_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   test UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
