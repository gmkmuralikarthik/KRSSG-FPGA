`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:07:25 12/11/2018 
// Design Name: 
// Module Name:    hallsensors 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module hallsencoders( hall,count,clk
    );

input clk,[2:0]hall,
output [7:0]count,

endmodule
